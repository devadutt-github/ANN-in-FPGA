module ann_tb;

  reg [19:0] img_tb[0:783];
  wire [9:0] out_tb[0:9];

  // Instantiate the design under test (DUT)
  ann dut (
    .img(img_tb),
    .out(out_tb)
  );

  // Provide initial values for img
 initial begin
img_tb[0] = 0 ;
img_tb[1] = 0 ;
img_tb[2] = 0 ;
img_tb[3] = 0 ;
img_tb[4] = 0 ;
img_tb[5] = 0 ;
img_tb[6] = 0 ;
img_tb[7] = 0 ;
img_tb[8] = 0 ;
img_tb[9] = 0 ;
img_tb[10] = 0 ;
img_tb[11] = 0 ;
img_tb[12] = 0 ;
img_tb[13] = 0 ;
img_tb[14] = 0 ;
img_tb[15] = 0 ;
img_tb[16] = 0 ;
img_tb[17] = 0 ;
img_tb[18] = 0 ;
img_tb[19] = 0 ;
img_tb[20] = 0 ;
img_tb[21] = 0 ;
img_tb[22] = 0 ;
img_tb[23] = 0 ;
img_tb[24] = 0 ;
img_tb[25] = 0 ;
img_tb[26] = 0 ;
img_tb[27] = 0 ;
img_tb[28] = 0 ;
img_tb[29] = 0 ;
img_tb[30] = 0 ;
img_tb[31] = 0 ;
img_tb[32] = 0 ;
img_tb[33] = 0 ;
img_tb[34] = 0 ;
img_tb[35] = 0 ;
img_tb[36] = 0 ;
img_tb[37] = 0 ;
img_tb[38] = 0 ;
img_tb[39] = 0 ;
img_tb[40] = 0 ;
img_tb[41] = 0 ;
img_tb[42] = 0 ;
img_tb[43] = 0 ;
img_tb[44] = 0 ;
img_tb[45] = 0 ;
img_tb[46] = 0 ;
img_tb[47] = 0 ;
img_tb[48] = 0 ;
img_tb[49] = 0 ;
img_tb[50] = 0 ;
img_tb[51] = 0 ;
img_tb[52] = 0 ;
img_tb[53] = 0 ;
img_tb[54] = 0 ;
img_tb[55] = 0 ;
img_tb[56] = 0 ;
img_tb[57] = 0 ;
img_tb[58] = 0 ;
img_tb[59] = 0 ;
img_tb[60] = 0 ;
img_tb[61] = 0 ;
img_tb[62] = 0 ;
img_tb[63] = 0 ;
img_tb[64] = 0 ;
img_tb[65] = 0 ;
img_tb[66] = 0 ;
img_tb[67] = 0 ;
img_tb[68] = 0 ;
img_tb[69] = 0 ;
img_tb[70] = 0 ;
img_tb[71] = 0 ;
img_tb[72] = 0 ;
img_tb[73] = 0 ;
img_tb[74] = 0 ;
img_tb[75] = 0 ;
img_tb[76] = 0 ;
img_tb[77] = 0 ;
img_tb[78] = 0 ;
img_tb[79] = 0 ;
img_tb[80] = 0 ;
img_tb[81] = 0 ;
img_tb[82] = 0 ;
img_tb[83] = 0 ;
img_tb[84] = 0 ;
img_tb[85] = 0 ;
img_tb[86] = 0 ;
img_tb[87] = 0 ;
img_tb[88] = 0 ;
img_tb[89] = 0 ;
img_tb[90] = 0 ;
img_tb[91] = 0 ;
img_tb[92] = 0 ;
img_tb[93] = 0 ;
img_tb[94] = 0 ;
img_tb[95] = 0 ;
img_tb[96] = 0 ;
img_tb[97] = 0 ;
img_tb[98] = 0 ;
img_tb[99] = 0 ;
img_tb[100] = 0 ;
img_tb[101] = 0 ;
img_tb[102] = 0 ;
img_tb[103] = 0 ;
img_tb[104] = 0 ;
img_tb[105] = 0 ;
img_tb[106] = 0 ;
img_tb[107] = 0 ;
img_tb[108] = 0 ;
img_tb[109] = 0 ;
img_tb[110] = 0 ;
img_tb[111] = 0 ;
img_tb[112] = 0 ;
img_tb[113] = 0 ;
img_tb[114] = 0 ;
img_tb[115] = 0 ;
img_tb[116] = 0 ;
img_tb[117] = 0 ;
img_tb[118] = 0 ;
img_tb[119] = 0 ;
img_tb[120] = 0 ;
img_tb[121] = 0 ;
img_tb[122] = 0 ;
img_tb[123] = 0 ;
img_tb[124] = 0 ;
img_tb[125] = 0 ;
img_tb[126] = 0 ;
img_tb[127] = 0 ;
img_tb[128] = 0 ;
img_tb[129] = 0 ;
img_tb[130] = 0 ;
img_tb[131] = 0 ;
img_tb[132] = 0 ;
img_tb[133] = 0 ;
img_tb[134] = 0 ;
img_tb[135] = 0 ;
img_tb[136] = 0 ;
img_tb[137] = 0 ;
img_tb[138] = 0 ;
img_tb[139] = 0 ;
img_tb[140] = 0 ;
img_tb[141] = 0 ;
img_tb[142] = 0 ;
img_tb[143] = 0 ;
img_tb[144] = 0 ;
img_tb[145] = 0 ;
img_tb[146] = 0 ;
img_tb[147] = 0 ;
img_tb[148] = 0 ;
img_tb[149] = 0 ;
img_tb[150] = 0 ;
img_tb[151] = 0 ;
img_tb[152] = 20 ;
img_tb[153] = 252 ;
img_tb[154] = 791 ;
img_tb[155] = 0 ;
img_tb[156] = 0 ;
img_tb[157] = 0 ;
img_tb[158] = 0 ;
img_tb[159] = 0 ;
img_tb[160] = 0 ;
img_tb[161] = 0 ;
img_tb[162] = 0 ;
img_tb[163] = 0 ;
img_tb[164] = 0 ;
img_tb[165] = 0 ;
img_tb[166] = 0 ;
img_tb[167] = 0 ;
img_tb[168] = 0 ;
img_tb[169] = 0 ;
img_tb[170] = 0 ;
img_tb[171] = 0 ;
img_tb[172] = 0 ;
img_tb[173] = 0 ;
img_tb[174] = 0 ;
img_tb[175] = 0 ;
img_tb[176] = 0 ;
img_tb[177] = 0 ;
img_tb[178] = 0 ;
img_tb[179] = 0 ;
img_tb[180] = 80 ;
img_tb[181] = 1019 ;
img_tb[182] = 923 ;
img_tb[183] = 96 ;
img_tb[184] = 0 ;
img_tb[185] = 0 ;
img_tb[186] = 0 ;
img_tb[187] = 0 ;
img_tb[188] = 0 ;
img_tb[189] = 0 ;
img_tb[190] = 0 ;
img_tb[191] = 0 ;
img_tb[192] = 0 ;
img_tb[193] = 0 ;
img_tb[194] = 0 ;
img_tb[195] = 0 ;
img_tb[196] = 0 ;
img_tb[197] = 0 ;
img_tb[198] = 0 ;
img_tb[199] = 0 ;
img_tb[200] = 0 ;
img_tb[201] = 0 ;
img_tb[202] = 0 ;
img_tb[203] = 0 ;
img_tb[204] = 0 ;
img_tb[205] = 0 ;
img_tb[206] = 0 ;
img_tb[207] = 0 ;
img_tb[208] = 80 ;
img_tb[209] = 1019 ;
img_tb[210] = 1019 ;
img_tb[211] = 192 ;
img_tb[212] = 0 ;
img_tb[213] = 0 ;
img_tb[214] = 0 ;
img_tb[215] = 0 ;
img_tb[216] = 0 ;
img_tb[217] = 0 ;
img_tb[218] = 0 ;
img_tb[219] = 0 ;
img_tb[220] = 0 ;
img_tb[221] = 0 ;
img_tb[222] = 0 ;
img_tb[223] = 0 ;
img_tb[224] = 0 ;
img_tb[225] = 0 ;
img_tb[226] = 0 ;
img_tb[227] = 0 ;
img_tb[228] = 0 ;
img_tb[229] = 0 ;
img_tb[230] = 0 ;
img_tb[231] = 0 ;
img_tb[232] = 0 ;
img_tb[233] = 0 ;
img_tb[234] = 0 ;
img_tb[235] = 0 ;
img_tb[236] = 80 ;
img_tb[237] = 1019 ;
img_tb[238] = 1024 ;
img_tb[239] = 192 ;
img_tb[240] = 0 ;
img_tb[241] = 0 ;
img_tb[242] = 0 ;
img_tb[243] = 0 ;
img_tb[244] = 0 ;
img_tb[245] = 0 ;
img_tb[246] = 0 ;
img_tb[247] = 0 ;
img_tb[248] = 0 ;
img_tb[249] = 0 ;
img_tb[250] = 0 ;
img_tb[251] = 0 ;
img_tb[252] = 0 ;
img_tb[253] = 0 ;
img_tb[254] = 0 ;
img_tb[255] = 0 ;
img_tb[256] = 0 ;
img_tb[257] = 0 ;
img_tb[258] = 0 ;
img_tb[259] = 0 ;
img_tb[260] = 0 ;
img_tb[261] = 0 ;
img_tb[262] = 0 ;
img_tb[263] = 0 ;
img_tb[264] = 80 ;
img_tb[265] = 1019 ;
img_tb[266] = 1019 ;
img_tb[267] = 228 ;
img_tb[268] = 0 ;
img_tb[269] = 0 ;
img_tb[270] = 0 ;
img_tb[271] = 0 ;
img_tb[272] = 0 ;
img_tb[273] = 0 ;
img_tb[274] = 0 ;
img_tb[275] = 0 ;
img_tb[276] = 0 ;
img_tb[277] = 0 ;
img_tb[278] = 0 ;
img_tb[279] = 0 ;
img_tb[280] = 0 ;
img_tb[281] = 0 ;
img_tb[282] = 0 ;
img_tb[283] = 0 ;
img_tb[284] = 0 ;
img_tb[285] = 0 ;
img_tb[286] = 0 ;
img_tb[287] = 0 ;
img_tb[288] = 0 ;
img_tb[289] = 0 ;
img_tb[290] = 0 ;
img_tb[291] = 0 ;
img_tb[292] = 80 ;
img_tb[293] = 1019 ;
img_tb[294] = 1019 ;
img_tb[295] = 433 ;
img_tb[296] = 0 ;
img_tb[297] = 0 ;
img_tb[298] = 0 ;
img_tb[299] = 0 ;
img_tb[300] = 0 ;
img_tb[301] = 0 ;
img_tb[302] = 0 ;
img_tb[303] = 0 ;
img_tb[304] = 0 ;
img_tb[305] = 0 ;
img_tb[306] = 0 ;
img_tb[307] = 0 ;
img_tb[308] = 0 ;
img_tb[309] = 0 ;
img_tb[310] = 0 ;
img_tb[311] = 0 ;
img_tb[312] = 0 ;
img_tb[313] = 0 ;
img_tb[314] = 0 ;
img_tb[315] = 0 ;
img_tb[316] = 0 ;
img_tb[317] = 0 ;
img_tb[318] = 0 ;
img_tb[319] = 0 ;
img_tb[320] = 64 ;
img_tb[321] = 959 ;
img_tb[322] = 1019 ;
img_tb[323] = 574 ;
img_tb[324] = 0 ;
img_tb[325] = 0 ;
img_tb[326] = 0 ;
img_tb[327] = 0 ;
img_tb[328] = 0 ;
img_tb[329] = 0 ;
img_tb[330] = 0 ;
img_tb[331] = 0 ;
img_tb[332] = 0 ;
img_tb[333] = 0 ;
img_tb[334] = 0 ;
img_tb[335] = 0 ;
img_tb[336] = 0 ;
img_tb[337] = 0 ;
img_tb[338] = 0 ;
img_tb[339] = 0 ;
img_tb[340] = 0 ;
img_tb[341] = 0 ;
img_tb[342] = 0 ;
img_tb[343] = 0 ;
img_tb[344] = 0 ;
img_tb[345] = 0 ;
img_tb[346] = 0 ;
img_tb[347] = 0 ;
img_tb[348] = 0 ;
img_tb[349] = 714 ;
img_tb[350] = 1019 ;
img_tb[351] = 574 ;
img_tb[352] = 0 ;
img_tb[353] = 0 ;
img_tb[354] = 0 ;
img_tb[355] = 0 ;
img_tb[356] = 0 ;
img_tb[357] = 0 ;
img_tb[358] = 0 ;
img_tb[359] = 0 ;
img_tb[360] = 0 ;
img_tb[361] = 0 ;
img_tb[362] = 0 ;
img_tb[363] = 0 ;
img_tb[364] = 0 ;
img_tb[365] = 0 ;
img_tb[366] = 0 ;
img_tb[367] = 0 ;
img_tb[368] = 0 ;
img_tb[369] = 0 ;
img_tb[370] = 0 ;
img_tb[371] = 0 ;
img_tb[372] = 0 ;
img_tb[373] = 0 ;
img_tb[374] = 0 ;
img_tb[375] = 0 ;
img_tb[376] = 0 ;
img_tb[377] = 714 ;
img_tb[378] = 1019 ;
img_tb[379] = 574 ;
img_tb[380] = 0 ;
img_tb[381] = 0 ;
img_tb[382] = 0 ;
img_tb[383] = 0 ;
img_tb[384] = 0 ;
img_tb[385] = 0 ;
img_tb[386] = 0 ;
img_tb[387] = 0 ;
img_tb[388] = 0 ;
img_tb[389] = 0 ;
img_tb[390] = 0 ;
img_tb[391] = 0 ;
img_tb[392] = 0 ;
img_tb[393] = 0 ;
img_tb[394] = 0 ;
img_tb[395] = 0 ;
img_tb[396] = 0 ;
img_tb[397] = 0 ;
img_tb[398] = 0 ;
img_tb[399] = 0 ;
img_tb[400] = 0 ;
img_tb[401] = 0 ;
img_tb[402] = 0 ;
img_tb[403] = 0 ;
img_tb[404] = 0 ;
img_tb[405] = 714 ;
img_tb[406] = 1019 ;
img_tb[407] = 650 ;
img_tb[408] = 0 ;
img_tb[409] = 0 ;
img_tb[410] = 0 ;
img_tb[411] = 0 ;
img_tb[412] = 0 ;
img_tb[413] = 0 ;
img_tb[414] = 0 ;
img_tb[415] = 0 ;
img_tb[416] = 0 ;
img_tb[417] = 0 ;
img_tb[418] = 0 ;
img_tb[419] = 0 ;
img_tb[420] = 0 ;
img_tb[421] = 0 ;
img_tb[422] = 0 ;
img_tb[423] = 0 ;
img_tb[424] = 0 ;
img_tb[425] = 0 ;
img_tb[426] = 0 ;
img_tb[427] = 0 ;
img_tb[428] = 0 ;
img_tb[429] = 0 ;
img_tb[430] = 0 ;
img_tb[431] = 0 ;
img_tb[432] = 0 ;
img_tb[433] = 714 ;
img_tb[434] = 1019 ;
img_tb[435] = 963 ;
img_tb[436] = 0 ;
img_tb[437] = 0 ;
img_tb[438] = 0 ;
img_tb[439] = 0 ;
img_tb[440] = 0 ;
img_tb[441] = 0 ;
img_tb[442] = 0 ;
img_tb[443] = 0 ;
img_tb[444] = 0 ;
img_tb[445] = 0 ;
img_tb[446] = 0 ;
img_tb[447] = 0 ;
img_tb[448] = 0 ;
img_tb[449] = 0 ;
img_tb[450] = 0 ;
img_tb[451] = 0 ;
img_tb[452] = 0 ;
img_tb[453] = 0 ;
img_tb[454] = 0 ;
img_tb[455] = 0 ;
img_tb[456] = 0 ;
img_tb[457] = 0 ;
img_tb[458] = 0 ;
img_tb[459] = 0 ;
img_tb[460] = 0 ;
img_tb[461] = 453 ;
img_tb[462] = 1019 ;
img_tb[463] = 963 ;
img_tb[464] = 0 ;
img_tb[465] = 0 ;
img_tb[466] = 0 ;
img_tb[467] = 0 ;
img_tb[468] = 0 ;
img_tb[469] = 0 ;
img_tb[470] = 0 ;
img_tb[471] = 0 ;
img_tb[472] = 0 ;
img_tb[473] = 0 ;
img_tb[474] = 0 ;
img_tb[475] = 0 ;
img_tb[476] = 0 ;
img_tb[477] = 0 ;
img_tb[478] = 0 ;
img_tb[479] = 0 ;
img_tb[480] = 0 ;
img_tb[481] = 0 ;
img_tb[482] = 0 ;
img_tb[483] = 0 ;
img_tb[484] = 0 ;
img_tb[485] = 0 ;
img_tb[486] = 0 ;
img_tb[487] = 0 ;
img_tb[488] = 0 ;
img_tb[489] = 333 ;
img_tb[490] = 1019 ;
img_tb[491] = 983 ;
img_tb[492] = 124 ;
img_tb[493] = 0 ;
img_tb[494] = 0 ;
img_tb[495] = 0 ;
img_tb[496] = 0 ;
img_tb[497] = 0 ;
img_tb[498] = 0 ;
img_tb[499] = 0 ;
img_tb[500] = 0 ;
img_tb[501] = 0 ;
img_tb[502] = 0 ;
img_tb[503] = 0 ;
img_tb[504] = 0 ;
img_tb[505] = 0 ;
img_tb[506] = 0 ;
img_tb[507] = 0 ;
img_tb[508] = 0 ;
img_tb[509] = 0 ;
img_tb[510] = 0 ;
img_tb[511] = 0 ;
img_tb[512] = 0 ;
img_tb[513] = 0 ;
img_tb[514] = 0 ;
img_tb[515] = 0 ;
img_tb[516] = 0 ;
img_tb[517] = 317 ;
img_tb[518] = 1019 ;
img_tb[519] = 987 ;
img_tb[520] = 152 ;
img_tb[521] = 0 ;
img_tb[522] = 0 ;
img_tb[523] = 0 ;
img_tb[524] = 0 ;
img_tb[525] = 0 ;
img_tb[526] = 0 ;
img_tb[527] = 0 ;
img_tb[528] = 0 ;
img_tb[529] = 0 ;
img_tb[530] = 0 ;
img_tb[531] = 0 ;
img_tb[532] = 0 ;
img_tb[533] = 0 ;
img_tb[534] = 0 ;
img_tb[535] = 0 ;
img_tb[536] = 0 ;
img_tb[537] = 0 ;
img_tb[538] = 0 ;
img_tb[539] = 0 ;
img_tb[540] = 0 ;
img_tb[541] = 0 ;
img_tb[542] = 0 ;
img_tb[543] = 0 ;
img_tb[544] = 0 ;
img_tb[545] = 0 ;
img_tb[546] = 859 ;
img_tb[547] = 1019 ;
img_tb[548] = 602 ;
img_tb[549] = 0 ;
img_tb[550] = 0 ;
img_tb[551] = 0 ;
img_tb[552] = 0 ;
img_tb[553] = 0 ;
img_tb[554] = 0 ;
img_tb[555] = 0 ;
img_tb[556] = 0 ;
img_tb[557] = 0 ;
img_tb[558] = 0 ;
img_tb[559] = 0 ;
img_tb[560] = 0 ;
img_tb[561] = 0 ;
img_tb[562] = 0 ;
img_tb[563] = 0 ;
img_tb[564] = 0 ;
img_tb[565] = 0 ;
img_tb[566] = 0 ;
img_tb[567] = 0 ;
img_tb[568] = 0 ;
img_tb[569] = 0 ;
img_tb[570] = 0 ;
img_tb[571] = 0 ;
img_tb[572] = 0 ;
img_tb[573] = 0 ;
img_tb[574] = 578 ;
img_tb[575] = 967 ;
img_tb[576] = 32 ;
img_tb[577] = 0 ;
img_tb[578] = 0 ;
img_tb[579] = 0 ;
img_tb[580] = 0 ;
img_tb[581] = 0 ;
img_tb[582] = 0 ;
img_tb[583] = 0 ;
img_tb[584] = 0 ;
img_tb[585] = 0 ;
img_tb[586] = 0 ;
img_tb[587] = 0 ;
img_tb[588] = 0 ;
img_tb[589] = 0 ;
img_tb[590] = 0 ;
img_tb[591] = 0 ;
img_tb[592] = 0 ;
img_tb[593] = 0 ;
img_tb[594] = 0 ;
img_tb[595] = 0 ;
img_tb[596] = 0 ;
img_tb[597] = 0 ;
img_tb[598] = 0 ;
img_tb[599] = 0 ;
img_tb[600] = 0 ;
img_tb[601] = 0 ;
img_tb[602] = 578 ;
img_tb[603] = 963 ;
img_tb[604] = 8 ;
img_tb[605] = 0 ;
img_tb[606] = 0 ;
img_tb[607] = 0 ;
img_tb[608] = 0 ;
img_tb[609] = 0 ;
img_tb[610] = 0 ;
img_tb[611] = 0 ;
img_tb[612] = 0 ;
img_tb[613] = 0 ;
img_tb[614] = 0 ;
img_tb[615] = 0 ;
img_tb[616] = 0 ;
img_tb[617] = 0 ;
img_tb[618] = 0 ;
img_tb[619] = 0 ;
img_tb[620] = 0 ;
img_tb[621] = 0 ;
img_tb[622] = 0 ;
img_tb[623] = 0 ;
img_tb[624] = 0 ;
img_tb[625] = 0 ;
img_tb[626] = 0 ;
img_tb[627] = 0 ;
img_tb[628] = 0 ;
img_tb[629] = 0 ;
img_tb[630] = 578 ;
img_tb[631] = 1019 ;
img_tb[632] = 329 ;
img_tb[633] = 0 ;
img_tb[634] = 0 ;
img_tb[635] = 0 ;
img_tb[636] = 0 ;
img_tb[637] = 0 ;
img_tb[638] = 0 ;
img_tb[639] = 0 ;
img_tb[640] = 0 ;
img_tb[641] = 0 ;
img_tb[642] = 0 ;
img_tb[643] = 0 ;
img_tb[644] = 0 ;
img_tb[645] = 0 ;
img_tb[646] = 0 ;
img_tb[647] = 0 ;
img_tb[648] = 0 ;
img_tb[649] = 0 ;
img_tb[650] = 0 ;
img_tb[651] = 0 ;
img_tb[652] = 0 ;
img_tb[653] = 0 ;
img_tb[654] = 0 ;
img_tb[655] = 0 ;
img_tb[656] = 0 ;
img_tb[657] = 0 ;
img_tb[658] = 923 ;
img_tb[659] = 991 ;
img_tb[660] = 160 ;
img_tb[661] = 0 ;
img_tb[662] = 0 ;
img_tb[663] = 0 ;
img_tb[664] = 0 ;
img_tb[665] = 0 ;
img_tb[666] = 0 ;
img_tb[667] = 0 ;
img_tb[668] = 0 ;
img_tb[669] = 0 ;
img_tb[670] = 0 ;
img_tb[671] = 0 ;
img_tb[672] = 0 ;
img_tb[673] = 0 ;
img_tb[674] = 0 ;
img_tb[675] = 0 ;
img_tb[676] = 0 ;
img_tb[677] = 0 ;
img_tb[678] = 0 ;
img_tb[679] = 0 ;
img_tb[680] = 0 ;
img_tb[681] = 0 ;
img_tb[682] = 0 ;
img_tb[683] = 0 ;
img_tb[684] = 0 ;
img_tb[685] = 0 ;
img_tb[686] = 674 ;
img_tb[687] = 839 ;
img_tb[688] = 124 ;
img_tb[689] = 0 ;
img_tb[690] = 0 ;
img_tb[691] = 0 ;
img_tb[692] = 0 ;
img_tb[693] = 0 ;
img_tb[694] = 0 ;
img_tb[695] = 0 ;
img_tb[696] = 0 ;
img_tb[697] = 0 ;
img_tb[698] = 0 ;
img_tb[699] = 0 ;
img_tb[700] = 0 ;
img_tb[701] = 0 ;
img_tb[702] = 0 ;
img_tb[703] = 0 ;
img_tb[704] = 0 ;
img_tb[705] = 0 ;
img_tb[706] = 0 ;
img_tb[707] = 0 ;
img_tb[708] = 0 ;
img_tb[709] = 0 ;
img_tb[710] = 0 ;
img_tb[711] = 0 ;
img_tb[712] = 0 ;
img_tb[713] = 0 ;
img_tb[714] = 0 ;
img_tb[715] = 0 ;
img_tb[716] = 0 ;
img_tb[717] = 0 ;
img_tb[718] = 0 ;
img_tb[719] = 0 ;
img_tb[720] = 0 ;
img_tb[721] = 0 ;
img_tb[722] = 0 ;
img_tb[723] = 0 ;
img_tb[724] = 0 ;
img_tb[725] = 0 ;
img_tb[726] = 0 ;
img_tb[727] = 0 ;
img_tb[728] = 0 ;
img_tb[729] = 0 ;
img_tb[730] = 0 ;
img_tb[731] = 0 ;
img_tb[732] = 0 ;
img_tb[733] = 0 ;
img_tb[734] = 0 ;
img_tb[735] = 0 ;
img_tb[736] = 0 ;
img_tb[737] = 0 ;
img_tb[738] = 0 ;
img_tb[739] = 0 ;
img_tb[740] = 0 ;
img_tb[741] = 0 ;
img_tb[742] = 0 ;
img_tb[743] = 0 ;
img_tb[744] = 0 ;
img_tb[745] = 0 ;
img_tb[746] = 0 ;
img_tb[747] = 0 ;
img_tb[748] = 0 ;
img_tb[749] = 0 ;
img_tb[750] = 0 ;
img_tb[751] = 0 ;
img_tb[752] = 0 ;
img_tb[753] = 0 ;
img_tb[754] = 0 ;
img_tb[755] = 0 ;
img_tb[756] = 0 ;
img_tb[757] = 0 ;
img_tb[758] = 0 ;
img_tb[759] = 0 ;
img_tb[760] = 0 ;
img_tb[761] = 0 ;
img_tb[762] = 0 ;
img_tb[763] = 0 ;
img_tb[764] = 0 ;
img_tb[765] = 0 ;
img_tb[766] = 0 ;
img_tb[767] = 0 ;
img_tb[768] = 0 ;
img_tb[769] = 0 ;
img_tb[770] = 0 ;
img_tb[771] = 0 ;
img_tb[772] = 0 ;
img_tb[773] = 0 ;
img_tb[774] = 0 ;
img_tb[775] = 0 ;
img_tb[776] = 0 ;
img_tb[777] = 0 ;
img_tb[778] = 0 ;
img_tb[779] = 0 ;
img_tb[780] = 0 ;
img_tb[781] = 0 ;
img_tb[782] = 0 ;
img_tb[783] = 0 ;

end


endmodule
